.WIDTH out=100
* Nodes 4-5 correspond to output4 (see gate at 116,-110)
* Nodes 6-7 correspond to 54 (see gate at 118,-92)
* Nodes 8-9 correspond to 92 (see gate at 119,-12)
* Nodes 10-11 correspond to 118 (see gate at 11,-44)
* Nodes 12-13 correspond to 64 (see gate at 32,-28)
* Nodes 14-15 correspond to 28 (see gate at 34,-90)
* Nodes 16-17 correspond to 7 (see gate at 40,-110)
* Nodes 18-19 correspond to input2 (see drain at 40,-120)

C1 11 0 0.073pf
C2 9 0 0.075pf
C3 5 0 0.052pf
C4 15 0 0.074pf
C5 13 0 0.068pf
M1 0 7 5 2 e l=4.0u w=16.0u
M2 1 5 5 2 d l=8.0u w=4.0u
M3 7 1 9 2 e l=4.0u w=4.0u
M4 9 9 1 2 d l=9.0u w=4.0u
M5 9 11 0 2 e l=4.0u w=8.0u
M6 11 13 0 2 e l=4.0u w=8.0u
M7 11 11 1 2 d l=9.0u w=4.0u
M8 1 13 13 2 d l=4.0u w=4.0u
M9 13 15 0 2 e l=4.0u w=16.0u
M10 15 17 0 2 e l=4.0u w=32.0u
M11 15 15 1 2 d l=4.0u w=4.0u
M12 19 1 17 2 e l=4.0u w=4.0u

* Initial conditions:
.ic v(17)=0
.ic v(11)=5
.ic v(7)=0
.ic v(9)=0
.ic v(5)=5
.ic v(15)=5
.ic v(13)=0
.ic v(19)=0

vin 19 0 pulse(0 5 0ns 0ns 0ns)
.tran .1ns 20ns
.print tran V(17) V(15) V(13) V(11) V(7) V(5) (0,5)
.end
