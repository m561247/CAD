STEPS deck from "bob:symbolic:contents;"
.options gmin=1p reltol=1m abstol=1p vntol=1u 
.options trtol=7 chgtol=10f pivtol=100f pivrel=1m 
.options numdgt=4 tnom=27 
.options itl1=100 itl2=50 itl4=10 cptime=0 
.options method=trapezoidal maxord=2 
.options defl=100u defw=100u defad=0 defas=0 
.model m3006 pmos VTO=-0.8 KP=3e-05
mi0 supply in out 1 m3006 W=4u L=2u 
+ AD=8p AS=8p PD=8u PS=8u 
.model m3043 nmos VTO=0.8 KP=7e-05
mi1 out in n0 0 m3043 W=4u L=2u 
+ AD=8p AS=8p PD=8u PS=8u 
CPn0 n0 0 24.4fFarad
CPsupply supply 0 21.4fFarad
CPin in 0 6.35fFarad
CPout out 0 47.5fFarad
*** cross cap n0 supply 0 --- small
*** cross cap n0 in 0 --- small
*** cross cap n0 out 0 --- small
*** cross cap supply in 0 --- small
*** cross cap supply out 0 --- small
*** cross cap in out 0 --- small
* Term Vdd   ( INPUT,SUPPLY) is node supply
vdd supply 0
+ DC 1.5 
* Term GND   ( INPUT,GROUND) is node n0
* Term in    ( INPUT,SIGNAL) is node in
?no_device_name? in 0
+ PWL(0 0  2n 1.5 4n 1.5 6n 0  )

* Term out   (OUTPUT,SIGNAL) is node out
.plot dc v(out)
.op
.tran 1n 10u 0 0.1n 


.plot tran in out

.end
