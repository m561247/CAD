STEPS input deck from example:schematic

vcc 1 0 dc 5
r0 1 2 330
r1 1 3 330

.model m635 npn IS=1e-16 BF=100 VA=33
q2 2 4 5 m635 1
q3 3 0 5 m635 1
r4 5 0 2100
v5 4 0 dc 2 

.width in = 3000
.width out = 80
.end
