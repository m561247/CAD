STEPS deck from "nand:symbolic:contents;"
.options gmin=1p reltol=1m abstol=1p vntol=1u 
.options trtol=7 chgtol=10f pivtol=0.1p pivrel=1m 
.options numdgt=4 tnom=27 
.options itl1=100 itl2=50 itl4=10 cptime=0 
.options method=trapezoidal maxord=2 
.options defl=0.1m defw=0.1m defad=0 defas=0 
** ERROR: Can't open user file ~/foo.spice
m0 out a supply supply pmos W=4u L=2u 
+ AD=8p AS=8p PD=4u PS=4u NRD=0.5 NRS=0.5 
mi2 n1 a 0 0 nmos W=4u L=2u 
+ AD=8p AS=8p PD=4u PS=4u NRD=0.5 NRS=0.5 
mi3 n1 b out 0 nmos W=4u L=2u 
+ AD=8p AS=8p PD=4u PS=4u NRD=0.5 NRS=0.5 
mi1 supply b out supply pmos W=4u L=2u 
+ AD=8p AS=8p PD=4u PS=4u NRD=0.5 NRS=0.5 
CPout out 0 47.8fFarad
*** cross cap a b 0.0889f --- small
*** cross cap a n1 0 --- small
*** cross cap a out 0.723f --- small
*** cross cap b n1 0 --- small
*** cross cap b out 0.723f --- small
*** cross cap n1 out 0 --- small
* Term Vdd   ( INPUT,SUPPLY) is node supply
vdd supply 0
+ DC 5 
* Term GND   ( INPUT,GROUND) is node  0
* Term out   (OUTPUT,SIGNAL) is node out
* Term a     ( INPUT,SIGNAL) is node  a
va a 0
+ DC 5 
+ PULSE(0 5 0 0 0 0.1u  0.2u) 

* Term b     ( INPUT,SIGNAL) is node  b
vb b 0
+ DC 0 
+ PULSE(0 5 0 0 0 50n  0.1u) 

** START MODELS
.model npn npn IS=1e-16 BF=100 VA=33
.model pnp pnp IS=1e-16 BF=100 VA=34
.model nmos nmos VTO=0.8 KP=7e-05
.model pmos pmos VTO=-0.8 KP=3e-05
.model diode D IS=1e-16
.model njfet njf VTO=2
.model pjfet pjf VTO=-2
** END MODELS
.op
.dc va 0 5 0.1 
.tran 1n 0.2u 0 1n 


.print tran a b out

.end
