* Nodes 4-5 correspond to Out (see gate at 1,1)
* Nodes 6-7 correspond to E (see gate at 1,1)
* Nodes 8-9 correspond to D (see gate at 1,1)
* Nodes 10-11 correspond to C (see gate at 1,1)
* Nodes 12-13 correspond to B (see gate at 1,1)
* Nodes 14-15 correspond to A (see gate at 1,1)
* Nodes 16-17 correspond to In (see gate at 1,1)

C1 5 0 .00001pf
M1 1 5 5 2 d l=16.0u w=4.0u
M2 0 7 5 2 e l=4.0u w=4.0u
M3 0 9 7 2 e l=4.0u w=4.0u
M4 1 7 7 2 d l=16.0u w=4.0u
M5 1 9 9 2 d l=16.0u w=4.0u
M6 0 11 9 2 e l=4.0u w=4.0u
M7 0 13 11 2 e l=4.0u w=4.0u
M8 1 11 11 2 d l=16.0u w=4.0u
M9 1 13 13 2 d l=16.0u w=4.0u
M10 0 15 13 2 e l=4.0u w=4.0u
M11 0 17 15 2 e l=4.0u w=4.0u
M12 1 15 15 2 d l=16.0u w=4.0u

* Initial conditions:
.ic v(15)=5.000000
.ic v(13)=0.000000
.ic v(11)=5.000000
.ic v(9)=0.000000
.ic v(7)=5.000000
.ic v(17)=0.000000
.ic v(5)=0.000000

vin 17 0 pulse(0 5 0ns 0ns 0ns)
.tran 0.05ns 10ns
.plot tran V(5) (0,5)
.end
