.WIDTH out=120
* Nodes 4-5 correspond to Out (see gate at 1,1)
* Nodes 6-7 correspond to E2 (see gate at 1,1)
* Nodes 8-9 correspond to E (see gate at 1,1)
* Nodes 10-11 correspond to D (see gate at 1,1)
* Nodes 12-13 correspond to C (see gate at 1,1)
* Nodes 14-15 correspond to B2 (see gate at 1,1)
* Nodes 16-17 correspond to B (see gate at 1,1)
* Nodes 18-19 correspond to A (see gate at 1,1)
* Nodes 20-21 correspond to In (see gate at 1,1)

C1 15 0 0.041pf
C2 19 0 0.990pf
C3 17 0 0.047pf
C4 13 0 0.040pf
C5 11 0 0.190pf
C6 9 0 0.047pf
C7 21 0 0.042pf
C8 7 0 0.041pf
C9 5 0 0.048pf
M1 1 5 5 2 d l=16.0u w=4.0u
M2 0 7 5 2 e l=4.0u w=4.0u
M3 7 1 9 2 e l=4.0u w=4.0u
M4 0 11 9 2 e l=4.0u w=4.0u
M5 1 9 9 2 d l=16.0u w=4.0u
M6 1 11 11 2 d l=16.0u w=4.0u
M7 0 13 11 2 e l=4.0u w=4.0u
M8 0 15 13 2 e l=4.0u w=4.0u
M9 1 13 13 2 d l=16.0u w=4.0u
M10 15 1 17 2 e l=4.0u w=4.0u
M11 1 17 17 2 d l=16.0u w=4.0u
M12 0 19 17 2 e l=4.0u w=4.0u
M13 0 21 19 2 e l=4.0u w=4.0u
M14 1 19 19 2 d l=16.0u w=4.0u

* Initial conditions:
.ic v(15)=0.000000
.ic v(19)=5.000000
.ic v(17)=0.000000
.ic v(13)=5.000000
.ic v(11)=0.000000
.ic v(9)=5.000000
.ic v(21)=0.000000
.ic v(7)=5.000000
.ic v(5)=0.000000

vin 21 0 pulse(0 5 0ns 0ns 0ns)
.tran 0.4ns 80ns
.print tran V(5) V(7) V(11) V(13) V(15) V(19) (0,5)
.end
