STEPS deck from "nor:symbolic:contents;"
mi2 0 a out 0 nmos W=6u L=2u 
+ AD=12p AS=12p PD=6u PS=6u NRD=0.333 NRS=0.333 
mi3 out b 0 0 nmos W=6u L=2u 
+ AD=12p AS=12p PD=6u PS=6u NRD=0.333 NRS=0.333 
mi1 n0 b out Vdd pmos W=12u L=2u 
+ AD=24p AS=24p PD=12u PS=12u NRD=0.166 NRS=0.166 
mi0 Vdd a n0 Vdd pmos W=12u L=2u 
+ AD=24p AS=24p PD=12u PS=12u NRD=0.166 NRS=0.166 
CPn0 n0 0 18fFarad
CPout out 0 0.175pFarad
CPa a 0 60.7fFarad
CPb b 0 77.6fFarad
* Term GND   ( INPUT,GROUND) is node  0
* Term Vdd   ( INPUT,SUPPLY) is node Vdd
Vdd Vdd 0
+ DC 5 
* Term a     ( INPUT,SIGNAL) is node  a
vaaa a 0
+ DC 5 
+ PULSE(0.1 4.9 0 0 0 50n  0.1u) 

* Term b     ( INPUT,SIGNAL) is node  b
vb b 0
+ DC 5 
+ PULSE(0 5 0 0 0 25n  50n) 

* Term out   (OUTPUT,SIGNAL) is node out
**** LOAD on formal terminal "out"
CLOADout out 0 100fFarad
RLOADout out 0 100kOhm

** START MODELS
.model npn npn IS=1e-16 BF=100 VA=33
.model pnp pnp IS=1e-16 BF=100 VA=34
.model nmos nmos VTO=0.8 KP=7e-05
.model pmos pmos VTO=-0.8 KP=3e-05
.model diode d IS=1e-16
.model njfet njf VTO=2
.model pjfet pjf VTO=-2
** END MODELS
.tran 1n 0.1u 0 0 


.print tran a b out

.end
